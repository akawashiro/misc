module pc (
    input logic clk,
    input logic [31:0] pc_in,
    output logic [31:0] pc_out
);
    always_ff @(posedge clk)
    begin
        pc_out <= pc_in;
    end
endmodule

module pc_plus_4 (
    input logic clk,
    input logic [31:0] pc_in,
    output logic [31:0] pc_out
);
    pc_out <= pc_in + 4;
endmodule
